`include "apb_config_db.sv"
`include "apb_tx.sv"
`include "apb_gen.sv"
`include "apb_bfm.sv"
`include "apb_mon.sv"
`include "apb_scb.sv"
`include "apb_env.sv"
`include "apb_test.sv"
`include "apb_intf.sv"
`include "apb_dut.sv"
`include "apb_tb_top.sv"
